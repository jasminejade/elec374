module con_ff_logic(input [31:0] busout, input [3:0] IR);
	