`timescale 1ns/10ps

module inout_tb;
	reg PCout, MARin, IncPC, Zin;
	reg Zlowout, PCin, Read, MDRin;
	reg MDRout, IRin;
	reg GRA, Rin;
	reg GRB, GRC, Inportout;
	reg clk, clr;
	reg RAM_read, RAM_write;
	reg [4:0] opcode;
	
	parameter Default = 4'b0000, T0 = 4'b0001, T1 = 4'b0010, T2 = 4'b0011, T3 = 4'b0100;
	reg [3:0] Present_state = Default;

datapath DUT(
	.PCout (PCout),
	.Zlowout (Zlowout),
	.MDRout (MDRout),
	.MARin (MARin),
	.Zin (Zin),
	.PCin (PCin),
	.MDRin (MDRin),
	.IRin (IRin),
	.IncPC (IncPC),
	.Read (Read),
	.clk (clk),
	.clr (clr),
	.RAM_read (RAM_read),
	.RAM_write (RAM_write),
	.opcode (opcode),
	.GRA (GRA),
	.GRB (GRB),
	.GRC (GRC),
	.Rin_logic (Rin),
	.INPORTout (Inportout)
);

// add test logic here
initial begin
	clr = 0;
	clk = 0;
	forever #10 clk = ~ clk;
end

always @(posedge clk) // finite state machine; if clock rising-edge
	begin
		case (Present_state)
			Default : #40 Present_state = T0;
			T0 : #40 Present_state = T1;
			T1 : #40 Present_state = T2;
			T2 : #40 Present_state = T3;
		endcase
	end
	
always @(Present_state) // do the required job in each state
	begin
		case (Present_state) // assert the required signals in each clock cycle
			Default: begin
				PCout <= 0; Zlowout <= 0; MDRout <= 0; // initialize the signals
				MARin <= 0; Zin <= 0; PCin <= 0; MDRin <= 0; IRin <= 0;
				IncPC <= 0; Read <= 0; opcode <= 0; RAM_read <= 0; RAM_write <= 0;
				GRA <= 0; GRB <= 0; Rin <= 0; GRC <= 0; Inportout <= 0;
			end
			T0: begin // see if you need to de-assert these signals
				#10 PCout <= 1; MARin <= 1; IncPC <= 1; Zin <= 1;
				#10 PCout <= 0; MARin <= 0; IncPC <= 0; Zin <= 0;
			end
			T1: begin
				#10 Zlowout <= 1; PCin <= 1; Read <= 1; RAM_read <= 1; MDRin <= 1; 
				// Mdatain = opcode for “ldi R1, $75”	
				#10 Zlowout <= 0; PCin <= 0; Read <= 0; RAM_read <= 0; MDRin <= 0; 
			end
			T2: begin
				#10 MDRout <= 1; IRin <= 1;
				#10 MDRout <= 0; IRin <= 0;
			end
			T3: begin
				#10 Inportout <= 1; GRA <= 1; Rin <= 1;
				#10 Inportout <= 0; GRA <= 0; Rin <= 0;
			end
		endcase
	end
endmodule 