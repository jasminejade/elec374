module rotate(
	input wire [31:0]		A, B,
	input wire				op,
	output wire [63:0]	Z
);
	reg [63:0] result;
	wire [4:0] N;
	assign N = B%32;
		
	always @(*) begin
		case(op)
			0 : result = (N == 31) ? {A[0:0], A[31:1]} : 
							 (N == 30) ? {A[1:0], A[31:2]} : 
							 (N == 29) ? {A[2:0], A[31:3]} : 
							 (N == 28) ? {A[3:0], A[31:4]} : 
							 (N == 27) ? {A[4:0], A[31:5]} : 
							 (N == 26) ? {A[5:0], A[31:6]} : 
							 (N == 25) ? {A[6:0], A[31:7]} : 
							 (N == 24) ? {A[7:0], A[31:8]} : 
							 (N == 23) ? {A[8:0], A[31:9]} : 
							 (N == 22) ? {A[9:0], A[31:10]} : 
							 (N == 21) ? {A[10:0], A[31:11]} : 
							 (N == 20) ? {A[11:0], A[31:12]} : 
							 (N == 19) ? {A[12:0], A[31:13]} : 
							 (N == 18) ? {A[13:0], A[31:14]} : 
							 (N == 17) ? {A[14:0], A[31:15]} : 
							 (N == 16) ? {A[15:0], A[31:16]} : 
							 (N == 15) ? {A[16:0], A[31:17]} : 
							 (N == 14) ? {A[17:0], A[31:18]} : 
							 (N == 13) ? {A[18:0], A[31:19]} : 
							 (N == 12) ? {A[19:0], A[31:20]} : 
							 (N == 11) ? {A[20:0], A[31:21]} : 
							 (N == 10) ? {A[21:0], A[31:22]} : 
							 (N == 9) ? {A[22:0], A[31:23]} : 
							 (N == 8) ? {A[23:0], A[31:24]} : 
							 (N == 7) ? {A[24:0], A[31:25]} : 
							 (N == 6) ? {A[25:0], A[31:26]} : 
							 (N == 5) ? {A[26:0], A[31:27]} : 
							 (N == 4) ? {A[27:0], A[31:28]} : 
							 (N == 3) ? {A[28:0], A[31:29]} : 
							 (N == 2) ? {A[29:0], A[31:30]} : 
							 (N == 1) ? {A[30:0], A[31:31]} : A;

			1 : result = (N == 31) ? {A[30:0], A[31:31]} :
							 (N == 30) ? {A[29:0], A[31:30]} : 
							 (N == 29) ? {A[28:0], A[31:29]} : 
							 (N == 28) ? {A[27:0], A[31:28]} : 
							 (N == 27) ? {A[26:0], A[31:27]} : 
							 (N == 26) ? {A[25:0], A[31:26]} : 
							 (N == 25) ? {A[24:0], A[31:25]} : 
							 (N == 24) ? {A[23:0], A[31:24]} : 
							 (N == 23) ? {A[22:0], A[31:23]} : 
							 (N == 22) ? {A[21:0], A[31:22]} : 
							 (N == 21) ? {A[20:0], A[31:21]} : 
							 (N == 20) ? {A[19:0], A[31:20]} : 
							 (N == 19) ? {A[18:0], A[31:19]} : 
							 (N == 18) ? {A[17:0], A[31:18]} : 
							 (N == 17) ? {A[16:0], A[31:17]} : 
							 (N == 16) ? {A[15:0], A[31:16]} : 
							 (N == 15) ? {A[14:0], A[31:15]} : 
							 (N == 14) ? {A[13:0], A[31:14]} : 
							 (N == 13) ? {A[12:0], A[31:13]} : 
							 (N == 12) ? {A[11:0], A[31:12]} : 
							 (N == 11) ? {A[10:0], A[31:11]} : 
							 (N == 10) ? {A[9:0], A[31:10]} : 
							 (N == 9) ? {A[8:0], A[31:9]} : 
							 (N == 8) ? {A[7:0], A[31:8]} : 
							 (N == 7) ? {A[6:0], A[31:7]} : 
							 (N == 6) ? {A[5:0], A[31:6]} : 
							 (N == 5) ? {A[4:0], A[31:5]} : 
							 (N == 4) ? {A[3:0], A[31:4]} : 
							 (N == 3) ? {A[2:0], A[31:3]} : 
							 (N == 2) ? {A[1:0], A[31:2]} : 
							 (N == 1) ? {A[0:0], A[31:1]} : A;
		endcase
	end
	assign Z = result;
endmodule
